module hs(a, b, diff, borrow); 
input a, b; 
output diff, borrow; 
xor (diff, a, b); 
and (borrow, ~a, b); 
endmodule 